module rx;

endmodule